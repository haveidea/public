module conf_dummy(
   output reg [7:0]                  owam_byte5,
   output reg [7:0]                  owam_byte6,
   output reg [7:0]                  owam_byte7,
   output reg onewire_crok,
   output reg onewire_ctok,
   output reg onewire_reok,
   output reg onewire_ppm,
   output reg [15:0] onewire_temp,
   output reg [15:0] onewire_ttrim
);

endmodule

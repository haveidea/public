`define    CLK2M4PERIOD    416   //ns
`define    CLK2M4RATIO     1
`define    CLK2M4DUTY      50
`define    CLK300PERIOD    3328  //ns
`define    CLK300RATIO     1
`define    CLK300DUTY      50
`define    PRESENCEMIN     60    //us
`define    PRESENCEMAX     240   //us
`define    CELSIUS0DEG     8'h00 //Celsius degree

